module top_module();
    initial begin
        $display("Hello, world!");
    end
endmodule